// Copyright (c) 2019 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// Authors:
// - Wolfgang Roenninger <wroennin@iis.ee.ethz.ch>
// - Andreas Kurth <akurth@iis.ee.ethz.ch>
// - Florian Zaruba <zarubaf@iis.ee.ethz.ch>

/// axi_xbar: Fully-connected AXI4+ATOP crossbar with an arbitrary number of slave and master ports.
/// See `doc/axi_xbar.md` for the documentation, including the definition of parameters and ports.
module axi_xbar
  import cf_math_pkg::idx_width;
#(
  /// Configuration struct for the crossbar see `axi_pkg` for fields and definitions.
  parameter axi_pkg::xbar_cfg_t Cfg = '0,
  /// Enable atomic operations support.
  parameter bit ATOPs = 1'b1,
  /// Connectivity matrix
  parameter bit [Cfg.NoSlvPorts-1:0][Cfg.NoMstPorts-1:0] Connectivity = '1,
  /// AXI4+ATOP AW channel struct type for the slave ports.
  parameter type slv_aw_chan_t = logic,
  /// AXI4+ATOP AW channel struct type for the master ports.
  parameter type mst_aw_chan_t = logic,
  /// AXI4+ATOP W channel struct type for all ports.
  parameter type w_chan_t = logic,
  /// AXI4+ATOP B channel struct type for the slave ports.
  parameter type slv_b_chan_t = logic,
  /// AXI4+ATOP B channel struct type for the master ports.
  parameter type mst_b_chan_t = logic,
  /// AXI4+ATOP AR channel struct type for the slave ports.
  parameter type slv_ar_chan_t = logic,
  /// AXI4+ATOP AR channel struct type for the master ports.
  parameter type mst_ar_chan_t = logic,
  /// AXI4+ATOP R channel struct type for the slave ports.
  parameter type slv_r_chan_t = logic,
  /// AXI4+ATOP R channel struct type for the master ports.
  parameter type mst_r_chan_t = logic,
  /// AXI4+ATOP request struct type for the slave ports.
  parameter type slv_req_t = logic,
  /// AXI4+ATOP response struct type for the slave ports.
  parameter type slv_resp_t = logic,
  /// AXI4+ATOP request struct type for the master ports.
  parameter type mst_req_t = logic,
  /// AXI4+ATOP response struct type for the master ports
  parameter type mst_resp_t = logic,
  /// Address rule type for the address decoders from `common_cells:addr_decode`.
  /// Example types are provided in `axi_pkg`.
  /// Required struct fields:
  /// ```
  /// typedef struct packed {
  ///   int unsigned idx;
  ///   axi_addr_t   start_addr;
  ///   axi_addr_t   end_addr;
  /// } rule_t;
  /// ```
  parameter type rule_t = axi_pkg::xbar_rule_64_t,
  localparam int unsigned MstPortsIdxWidth = (Cfg.NoMstPorts == 32'd1) ? 32'd1 : unsigned'($clog2(
      Cfg.NoMstPorts
  ))
) (
  /// Clock, positive edge triggered.
  input  logic                                                  clk_i,
  /// Asynchronous reset, active low.
  input  logic                                                  rst_ni,
  /// Testmode enable, active high.
  input  logic                                                  test_i,
  /// AXI4+ATOP requests to the slave ports.
  input  slv_req_t  [ Cfg.NoSlvPorts-1:0]                       slv_ports_req_i,
  /// AXI4+ATOP responses of the slave ports.
  output slv_resp_t [ Cfg.NoSlvPorts-1:0]                       slv_ports_resp_o,
  /// AXI4+ATOP requests of the master ports.
  output mst_req_t  [ Cfg.NoMstPorts-1:0]                       mst_ports_req_o,
  /// AXI4+ATOP responses to the master ports.
  input  mst_resp_t [ Cfg.NoMstPorts-1:0]                       mst_ports_resp_i,
  /// Address map array input for the crossbar. This map is global for the whole module.
  /// It is used for routing the transactions to the respective master ports.
  /// Each master port can have multiple different rules.
  input  rule_t     [Cfg.NoAddrRules-1:0]                       addr_map_i,
  /// Enable default master port.
  input  logic      [ Cfg.NoSlvPorts-1:0]                       en_default_mst_port_i,
  /// Enables a default master port for each slave port. When this is enabled unmapped
  /// transactions get issued at the master port given by `default_mst_port_i`.
  /// When not used, tie to `'0`.
  input  logic      [ Cfg.NoSlvPorts-1:0][MstPortsIdxWidth-1:0] default_mst_port_i
);

  // signals into the axi_muxes, are of type slave as the multiplexer extends the ID
  slv_req_t  [Cfg.NoMstPorts-1:0][Cfg.NoSlvPorts-1:0] mst_reqs;
  slv_resp_t [Cfg.NoMstPorts-1:0][Cfg.NoSlvPorts-1:0] mst_resps;

  axi_xbar_unmuxed #(
    .Cfg         (Cfg),
    .ATOPs       (ATOPs),
    .Connectivity(Connectivity),
    .aw_chan_t   (slv_aw_chan_t),
    .w_chan_t    (w_chan_t),
    .b_chan_t    (slv_b_chan_t),
    .ar_chan_t   (slv_ar_chan_t),
    .r_chan_t    (slv_r_chan_t),
    .req_t       (slv_req_t),
    .resp_t      (slv_resp_t),
    .rule_t      (rule_t)
  ) i_xbar_unmuxed (
    .clk_i,
    .rst_ni,
    .test_i,
    .slv_ports_req_i,
    .slv_ports_resp_o,
    .mst_ports_req_o (mst_reqs),
    .mst_ports_resp_i(mst_resps),
    .addr_map_i,
    .en_default_mst_port_i,
    .default_mst_port_i
  );

  for (genvar i = 0; i < Cfg.NoMstPorts; i++) begin : gen_mst_port_mux
    axi_mux #(
      .SlvAxiIDWidth(Cfg.AxiIdWidthSlvPorts),  // ID width of the slave ports
      .slv_aw_chan_t(slv_aw_chan_t),           // AW Channel Type, slave ports
      .mst_aw_chan_t(mst_aw_chan_t),           // AW Channel Type, master port
      .w_chan_t     (w_chan_t),                //  W Channel Type, all ports
      .slv_b_chan_t (slv_b_chan_t),            //  B Channel Type, slave ports
      .mst_b_chan_t (mst_b_chan_t),            //  B Channel Type, master port
      .slv_ar_chan_t(slv_ar_chan_t),           // AR Channel Type, slave ports
      .mst_ar_chan_t(mst_ar_chan_t),           // AR Channel Type, master port
      .slv_r_chan_t (slv_r_chan_t),            //  R Channel Type, slave ports
      .mst_r_chan_t (mst_r_chan_t),            //  R Channel Type, master port
      .slv_req_t    (slv_req_t),
      .slv_resp_t   (slv_resp_t),
      .mst_req_t    (mst_req_t),
      .mst_resp_t   (mst_resp_t),
      .NoSlvPorts   (Cfg.NoSlvPorts),          // Number of Masters for the module
      .MaxWTrans    (Cfg.MaxSlvTrans),
      .FallThrough  (Cfg.FallThrough),
      .SpillAw      (Cfg.LatencyMode[4]),
      .SpillW       (Cfg.LatencyMode[3]),
      .SpillB       (Cfg.LatencyMode[2]),
      .SpillAr      (Cfg.LatencyMode[1]),
      .SpillR       (Cfg.LatencyMode[0])
    ) i_axi_mux (
      .clk_i,  // Clock
      .rst_ni,  // Asynchronous reset active low
      .test_i,  // Test Mode enable
      .slv_reqs_i (mst_reqs[i]),
      .slv_resps_o(mst_resps[i]),
      .mst_req_o  (mst_ports_req_o[i]),
      .mst_resp_i (mst_ports_resp_i[i])
    );
  end

  // pragma translate_off
`ifndef VERILATOR
`ifndef XSIM
  initial begin : check_params
    id_slv_req_ports :
    assert ($bits(slv_ports_req_i[0].aw.id) == Cfg.AxiIdWidthSlvPorts)
    else $fatal(1, $sformatf("Slv_req and aw_chan id width not equal."));
    id_slv_resp_ports :
    assert ($bits(slv_ports_resp_o[0].r.id) == Cfg.AxiIdWidthSlvPorts)
    else $fatal(1, $sformatf("Slv_req and aw_chan id width not equal."));
  end
`endif
`endif
  // pragma translate_on
endmodule

`include "axi/assign.svh"
`include "axi/typedef.svh"

module axi_xbar_intf
  import cf_math_pkg::idx_width;
#(
  parameter int unsigned AXI_USER_WIDTH = 0,
  parameter axi_pkg::xbar_cfg_t Cfg = '0,
  parameter bit ATOPS = 1'b1,
  parameter bit [Cfg.NoSlvPorts-1:0][Cfg.NoMstPorts-1:0] CONNECTIVITY = '1,
  parameter type rule_t = axi_pkg::xbar_rule_64_t,
  localparam int unsigned MstPortsIdxWidth = (Cfg.NoMstPorts == 32'd1) ? 32'd1 : unsigned'($clog2(
      Cfg.NoMstPorts
  ))
) (
  input logic clk_i,
  input logic rst_ni,
  input logic test_i,
  AXI_BUS.Slave slv_ports[Cfg.NoSlvPorts-1:0],
  AXI_BUS.Master mst_ports[Cfg.NoMstPorts-1:0],
  input rule_t [Cfg.NoAddrRules-1:0] addr_map_i,
  input logic [Cfg.NoSlvPorts-1:0] en_default_mst_port_i,
  input logic [Cfg.NoSlvPorts-1:0][MstPortsIdxWidth-1:0] default_mst_port_i
);

  localparam int unsigned AxiIdWidthMstPorts = Cfg.AxiIdWidthSlvPorts + $clog2(Cfg.NoSlvPorts);

  typedef logic [AxiIdWidthMstPorts     -1:0] id_mst_t;
  typedef logic [Cfg.AxiIdWidthSlvPorts -1:0] id_slv_t;
  typedef logic [Cfg.AxiAddrWidth       -1:0] addr_t;
  typedef logic [Cfg.AxiDataWidth       -1:0] data_t;
  typedef logic [Cfg.AxiDataWidth/8     -1:0] strb_t;
  typedef logic [AXI_USER_WIDTH         -1:0] user_t;

  `AXI_TYPEDEF_AW_CHAN_T(mst_aw_chan_t, addr_t, id_mst_t, user_t)
  `AXI_TYPEDEF_AW_CHAN_T(slv_aw_chan_t, addr_t, id_slv_t, user_t)
  `AXI_TYPEDEF_W_CHAN_T(w_chan_t, data_t, strb_t, user_t)
  `AXI_TYPEDEF_B_CHAN_T(mst_b_chan_t, id_mst_t, user_t)
  `AXI_TYPEDEF_B_CHAN_T(slv_b_chan_t, id_slv_t, user_t)
  `AXI_TYPEDEF_AR_CHAN_T(mst_ar_chan_t, addr_t, id_mst_t, user_t)
  `AXI_TYPEDEF_AR_CHAN_T(slv_ar_chan_t, addr_t, id_slv_t, user_t)
  `AXI_TYPEDEF_R_CHAN_T(mst_r_chan_t, data_t, id_mst_t, user_t)
  `AXI_TYPEDEF_R_CHAN_T(slv_r_chan_t, data_t, id_slv_t, user_t)
  `AXI_TYPEDEF_REQ_T(mst_req_t, mst_aw_chan_t, w_chan_t, mst_ar_chan_t)
  `AXI_TYPEDEF_REQ_T(slv_req_t, slv_aw_chan_t, w_chan_t, slv_ar_chan_t)
  `AXI_TYPEDEF_RESP_T(mst_resp_t, mst_b_chan_t, mst_r_chan_t)
  `AXI_TYPEDEF_RESP_T(slv_resp_t, slv_b_chan_t, slv_r_chan_t)

  mst_req_t  [Cfg.NoMstPorts-1:0] mst_reqs;
  mst_resp_t [Cfg.NoMstPorts-1:0] mst_resps;
  slv_req_t  [Cfg.NoSlvPorts-1:0] slv_reqs;
  slv_resp_t [Cfg.NoSlvPorts-1:0] slv_resps;

  for (genvar i = 0; i < Cfg.NoMstPorts; i++) begin : gen_assign_mst
    `AXI_ASSIGN_FROM_REQ(mst_ports[i], mst_reqs[i])
    `AXI_ASSIGN_TO_RESP(mst_resps[i], mst_ports[i])
  end

  for (genvar i = 0; i < Cfg.NoSlvPorts; i++) begin : gen_assign_slv
    `AXI_ASSIGN_TO_REQ(slv_reqs[i], slv_ports[i])
    `AXI_ASSIGN_FROM_RESP(slv_ports[i], slv_resps[i])
  end

  axi_xbar #(
    .Cfg          (Cfg),
    .ATOPs        (ATOPS),
    .Connectivity (CONNECTIVITY),
    .slv_aw_chan_t(slv_aw_chan_t),
    .mst_aw_chan_t(mst_aw_chan_t),
    .w_chan_t     (w_chan_t),
    .slv_b_chan_t (slv_b_chan_t),
    .mst_b_chan_t (mst_b_chan_t),
    .slv_ar_chan_t(slv_ar_chan_t),
    .mst_ar_chan_t(mst_ar_chan_t),
    .slv_r_chan_t (slv_r_chan_t),
    .mst_r_chan_t (mst_r_chan_t),
    .slv_req_t    (slv_req_t),
    .slv_resp_t   (slv_resp_t),
    .mst_req_t    (mst_req_t),
    .mst_resp_t   (mst_resp_t),
    .rule_t       (rule_t)
  ) i_xbar (
    .clk_i,
    .rst_ni,
    .test_i,
    .slv_ports_req_i (slv_reqs),
    .slv_ports_resp_o(slv_resps),
    .mst_ports_req_o (mst_reqs),
    .mst_ports_resp_i(mst_resps),
    .addr_map_i,
    .en_default_mst_port_i,
    .default_mst_port_i
  );

endmodule
